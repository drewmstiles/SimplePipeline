
module Adder(
	input [31:0] PCout,
	output reg[31:0] PCin
    );

	always @(PCout) begin

	end

endmodule
