module IM(
	input[31:0] PCout,
	output reg[31:0] IMout
    );

	reg [7:0] IM [0:39]; // 40 instructions, 1 word each, byte thin

	always @(PCout) begin
		assign IMout = {IM[PCout[31:0] + 0], IM[PCout[31:0] + 1], IM[PCout[31:0] + 2], IM[PCout[31:0] + 3]};
	end
	
	initial begin
	
IM[0] = 8'b10001100;
IM[1] = 8'b00000101;
IM[2] = 8'b00000000;
IM[3] = 8'b00000000;
IM[4] = 8'b10001100;
IM[5] = 8'b00001010;
IM[6] = 8'b00000000;
IM[7] = 8'b00000100;
IM[8] = 8'b00000000;
IM[9] = 8'b10101010;
IM[10] = 8'b01101000;
IM[11] = 8'b00100000;
IM[12] = 8'b10101100;
IM[13] = 8'b00001101;
IM[14] = 8'b00000000;
IM[15] = 8'b00001100;
IM[16] = 8'b00000000;
IM[17] = 8'b10101010;
IM[18] = 8'b01101000;
IM[19] = 8'b00100010;
IM[20] = 8'b10101100;
IM[21] = 8'b00001101;
IM[22] = 8'b00000000;
IM[23] = 8'b00010000;
IM[24] = 8'b00000000;
IM[25] = 8'b10101010;
IM[26] = 8'b01101000;
IM[27] = 8'b00100100;
IM[28] = 8'b10101100;
IM[29] = 8'b00001101;
IM[30] = 8'b00000000;
IM[31] = 8'b00010100;
IM[32] = 8'b00000000;
IM[33] = 8'b10101010;
IM[34] = 8'b01101000;
IM[35] = 8'b00100101;
IM[36] = 8'b10101100;
IM[37] = 8'b00001101;
IM[38] = 8'b00000000;
IM[39] = 8'b00011000;

	end
	
endmodule
